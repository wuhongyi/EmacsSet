// test.v --- 
// 
// Description: 
// Author: Hongyi Wu(吴鸿毅)
// Email: wuhongyi@qq.com 
// Created: 一 7月  2 03:17:27 2018 (+0800)
// Last-Updated: 一 7月  2 03:31:52 2018 (+0800)
//           By: Hongyi Wu(吴鸿毅)
//     Update #: 1
// URL: http://wuhongyi.cn 

module name
  (
   input clk;
   input rst_n;
   // output ;
   );
   
   // wire ;                  
   // reg ;

   // 连续赋值
   // assign  = ;
   
   // always 块
   
   // 模块h例化

endmodule

// 
// test.v ends here
